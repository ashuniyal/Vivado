`timescale 1ns / 1ps

module comp(input a,input b,output c);
xnor(c,a,b);
endmodule
